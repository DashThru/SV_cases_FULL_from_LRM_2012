////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        198
// Description: the continuous assignment statement 
// Note:        
//
////////////////////////////////////////////////////////////////



module adder (sum_out, carry_out, carry_in, ina, inb);
  output [3:0] sum_out;
  output carry_out;
  input [3:0] ina, inb;
  input carry_in;
  wire carry_out, carry_in;
  wire [3:0] sum_out, ina, inb;
  assign {carry_out, sum_out} = ina + inb + carry_in;
endmodule

module select_bus(busout, bus0, bus1, bus2, bus3, enable, s);
  parameter n = 16;
  parameter Zee = 16'bz;
  output [1:n] busout;
  input [1:n] bus0, bus1, bus2, bus3; input enable;
  input [1:2] s;
  tri [1:n] data; // net declaration
  // net declaration with continuous assignment
  tri [1:n] busout = enable ? data : Zee;
       // assignment statement with four continuous assignments
  assign
    data = (s == 0) ? bus0 : Zee,
    data = (s == 1) ? bus1 : Zee,
    data = (s == 2) ? bus2 : Zee,
    data = (s == 3) ? bus3 : Zee;
endmodule

module sv12_lrm_p0198_wire_mynet;
  wire mynet,enable;
  wire #10 wireA;
  assign (strong1, pull0) mynet = enable;

endmodule : sv12_lrm_p0198_wire_mynet
