////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        178
// Description: begin end blockb block name
// Note:        
//
////////////////////////////////////////////////////////////////

module sv12_lrm_p0178_begin_blockb_block;

  initial   
  begin: blockB // block name after the begin or fork ...
  end: blockB

endmodule : sv12_lrm_p0178_begin_blockb_block
