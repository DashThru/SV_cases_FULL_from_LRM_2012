////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        519
// Description: defining the coverage model: covergroup
// Note:        
//
////////////////////////////////////////////////////////////////

module sv12_lrm_p0519_covergroup_cg_endgroup;

  covergroup cg; endgroup
  cg cg_inst = new;

endmodule : sv12_lrm_p0519_covergroup_cg_endgroup
