////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        69
// Description: int unsigned ui
// Note:        
//
////////////////////////////////////////////////////////////////

module sv12_lrm_p0069_int_unsigned_ui;

  int unsigned ui;
  int signed si;
  
  chandle variable_name ;

endmodule : sv12_lrm_p0069_int_unsigned_ui
