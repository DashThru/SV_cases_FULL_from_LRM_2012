////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        12
// Description: program port declaration
// Note:        
//
////////////////////////////////////////////////////////////////

module sv12_lrm_p0012_program_test;
  // program instance
  sv12_lrm_p0012_program_test_p p_inst();
endmodule

program sv12_lrm_p0012_program_test_p (input clk, input [16:1] addr, inout [7:0] data);
  initial begin
  end
endprogram

