////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        233
// Description: shift operators
// Note:        
//
////////////////////////////////////////////////////////////////

module shift;
  logic [3:0] start, result;
  initial begin
    start = 1;
    result = (start << 2);
  end
endmodule

module ashift;
  logic signed [3:0] start, result;
  initial begin
    start = 4'b1000;
    result = (start >>> 2);
  end
endmodule

module sv12_lrm_p0233_module_shift;

  shift u_shift();
  ashift u_ashift();

endmodule : sv12_lrm_p0233_module_shift
