////////////////////////////////////////////////////////////////
//
// LRM:         SV2012
// Page:        446
// Description: expect statement and concurrent assertions
// Note:        
//
////////////////////////////////////////////////////////////////

program tst;
  logic clk,a,b,c;
  
  initial begin
    # 200ms;
    expect( @(posedge clk) a ##1 b ##1 c ) else $error( "expect failed" );
  end
endprogram

module A;
  logic a, clk;
  clocking cb_with_input @(posedge clk);
    input a;
    property p1;
	  a;
    endproperty
  endclocking
  clocking cb_without_input @(posedge clk);
    property p1;
      a;
    endproperty
  endclocking
  property p1;
    @(posedge clk) a;
  endproperty
  property p2;
    @(posedge clk) cb_with_input.a;
  endproperty
  a1: assert property (p1);
  a2: assert property (cb_with_input.p1);
  a3: assert property (p2);
  a4: assert property (cb_without_input.p1);
endmodule

module sv12_lrm_p0446_program_tst;

  logic clk;
  integer data;

  task automatic wait_for( integer value, output bit success );
  expect( @(posedge clk) ##[1:10] data == value ) success = 1;
    else success = 0;
  endtask
  initial begin
    bit ok;
    wait_for( 23, ok ); // wait for the value 23
  end

  A uA(); 

endmodule : sv12_lrm_p0446_program_tst
